/*MAS: 00 B  //  01 H  //  10 w  // 11 undefined
1 = read  //  0 = write
changed mem value for test purposes */

module ram512x8 (output reg [31:0]dataOut, output reg done, input enable, readWrite, input [8:0]address, input [31:0]dataIn, input [1:0]MAS);
	reg [8:0]mem[0:512];
	always @ (enable, readWrite, MAS, dataIn, address)
	begin
		if (enable)
		begin
			done = 0;
			if (readWrite) begin
				//Reading
				case(MAS)
<<<<<<< HEAD
					2'b00:	begin
						// case(address[1:0])
						// 	2'b00:	dataOut[7:0] = mem[address + 8'b0000011][7:0];
						// 	2'b01:	dataOut[7:0] = mem[address + 8'b0000010][7:0];
						// 	2'b10:	dataOut[7:0] = mem[address + 8'b0000001][7:0];
							//2'b11:	
							dataOut[7:0] = mem[address][7:0];
						//  endcase
=======
					2'b00:	begin // #15;
						case(A)
							2'b00:	dataOut[7:0] = mem[address + 8'b0000011][7:0];
							2'b01:	dataOut[7:0] = mem[address + 8'b0000010][7:0];
							2'b10:	dataOut[7:0] = mem[address + 8'b0000001][7:0];
							2'b11:	dataOut[7:0] = mem[address][7:0];
						endcase
>>>>>>> e5dd09604a2f15378edc301521c6fdc52121ca21
						dataOut[31:8] = 24'b0000_0000_0000_0000_0000_0000;
						
					end
<<<<<<< HEAD
					2'b01:	begin	
						// case(address[1])
						// 	1'b0:	begin
						// 		dataOut[15:8] = mem[address + 8'b0000010][7:0];
						// 		dataOut[7:0] = mem[address + 8'b0000011][7:0];
						// 	end
						// 	1'b1:	begin
=======
					2'b01:	begin // #20;
						case(A[1])
							1'b0:	begin
								dataOut[15:8] = mem[address + 8'b0000010][7:0];
								dataOut[7:0] = mem[address + 8'b0000011][7:0];
							end
							1'b1:	begin
>>>>>>> e5dd09604a2f15378edc301521c6fdc52121ca21
								dataOut[15:8] = mem[address][7:0];
								dataOut[7:0] = mem[address + 8'b0000001][7:0];
						//	end
						//endcase
						dataOut[31:16] = 16'b0000_0000_0000_0000;
						
					end
					2'b10:	begin // #30;
						dataOut[31:0] = {mem[address][7:0], 
										 mem[address + 8'b0000001][7:0], 
										 mem[address + 8'b0000010][7:0], 
										 mem[address + 8'b0000011][7:0]};
						
					end
					default: dataOut = dataOut;
				endcase
			end
			else begin
				//Writing
				case(MAS)
<<<<<<< HEAD
					2'b00:	begin	
						// case(A)
						// 	2'b00:	mem[address + 8'b0000011][7:0] = dataIn[7:0];
						// 	2'b01:	mem[address + 8'b0000010][7:0] = dataIn[7:0];
						// 	2'b10:	mem[address + 8'b0000001][7:0] = dataIn[7:0];
							// 2'b11:	
							mem[address][7:0] = dataIn[7:0];
						// endcase
						// #25;
					end
					2'b01:	begin
						// case(A[1])
						// 	1'b0:	begin
						// 		mem[address + 8'b0000010][7:0] = dataIn[15:8];
						// 		mem[address + 8'b0000011][7:0] = dataIn[7:0];
						// 	end
							// 1'b1:	begin
								mem[address][7:0] = dataIn[15:8];
								mem[address + 8'b0000001][7:0] = dataIn[7:0] ;
							// end
						// endcase
						//#35;
=======
					2'b00:	begin // #25;
						case(A)
							2'b00:	mem[address + 8'b0000011][7:0] = dataIn[7:0];
							2'b01:	mem[address + 8'b0000010][7:0] = dataIn[7:0];
							2'b10:	mem[address + 8'b0000001][7:0] = dataIn[7:0];
							2'b11:	mem[address][7:0] = dataIn[7:0];
						endcase
						
					end
					2'b01:	begin //#35;
						case(A[1])
							1'b0:	begin
								mem[address + 8'b0000010][7:0] = dataIn[15:8];
								mem[address + 8'b0000011][7:0] = dataIn[7:0];
							end
							1'b1:	begin
								mem[address][7:0] = dataIn[15:8];
								mem[address + 8'b0000001][7:0] = dataIn[7:0] ;
							end
						endcase
						
>>>>>>> e5dd09604a2f15378edc301521c6fdc52121ca21
					end
					2'b10:	begin //#60;
						mem[address + 8'b00000011][7:0] = dataIn[7:0];
						mem[address + 8'b00000010][7:0] = dataIn[15:8];
						mem[address + 8'b00000001][7:0] = dataIn[23:16];
						mem[address][7:0] = dataIn[31:24];
						
					end
					default: dataOut = dataOut;
				endcase
			end
			done = 1;
		end
		else
			dataOut = 32'bz;
	end
endmodule